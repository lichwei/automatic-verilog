    always@(*) begin
         
    end
