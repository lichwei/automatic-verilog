    always@(posedge clk or negedge rst_n) begin
        if(!rst_n)
             
        else 
             
    end
